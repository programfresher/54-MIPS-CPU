module INSTR(
input [31:0]instruction,
output [5:0]op,
output [4:0]rs,
output [4:0]rt,
output [4:0]rd,
output [4:0]shamt,
output [5:0]func,
output [15:0]imme16,
output [25:0]imme26
    );

assign op=instruction[31:26];
assign rs=instruction[25:21];
assign rt=instruction[20:16];
assign rd=instruction[15:11];
assign shamt=instruction[10:6];
assign func=instruction[5:0];
assign imme16=instruction[15:0];
assign imme26=instruction[25:0];

endmodule
